//contains all the sequence files including virtual sequence (named as p_seq)
package seq_pkg;

    import uvm_pkg::*;

    `include "uvm_macros.svh"

    `include "/home/abdullah_hassaan/Documents/Coverage_check_xbar_l2/Coverage_check_xbar_l2/xbar_latest1_coverage_extnd/xbar_latest/dv/seq_lib/seq_master.sv"
    
    `include "/home/abdullah_hassaan/Documents/Coverage_check_xbar_l2/Coverage_check_xbar_l2/xbar_latest1_coverage_extnd/xbar_latest/dv/seq_lib/seq_slave.sv"  
   
    `include "/home/abdullah_hassaan/Documents/Coverage_check_xbar_l2/Coverage_check_xbar_l2/xbar_latest1_coverage_extnd/xbar_latest/dv/seq_lib/p_seq.sv"
  
endpackage : seq_pkg
